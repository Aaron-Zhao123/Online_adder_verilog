library verilog;
use verilog.vl_types.all;
entity D_flipflop_with_initial is
    port(
        clk             : in     vl_logic;
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end D_flipflop_with_initial;
